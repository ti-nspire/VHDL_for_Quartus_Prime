library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.types.all;

entity coeffs_list is
	port(
		outp : out coefficient_array(0 to 100)(15 downto 0)
	);
end entity;

architecture rtl of coeffs_list is
begin
	outp <=
	
((16d"65519"),(16d"65524"),(16d"0"),(16d"14"),(16d"21"),(16d"17"),(16d"0"),(16d"65515"),(16d"65502"),(16d"65509"),(16d"0"),(16d"35"),(16d"56"),(16d"45"),(16d"0"),(16d"65479"),(16d"65446"),(16d"65465"),(16d"0"),(16d"88"),(16d"138"),(16d"108"),(16d"0"),(16d"65404"),(16d"65331"),(16d"65377"),(16d"0"),(16d"192"),(16d"297"),(16d"230"),(16d"0"),(16d"65261"),(16d"65109"),(16d"65205"),(16d"0"),(16d"399"),(16d"621"),(16d"485"),(16d"0"),(16d"64936"),(16d"64584"),(16d"64775"),(16d"0"),(16d"1008"),(16d"1683"),(16d"1443"),(16d"0"),(16d"63096"),(16d"60337"),(16d"58164"),(16d"24588"),(16d"58164"),(16d"60337"),(16d"63096"),(16d"0"),(16d"1443"),(16d"1683"),(16d"1008"),(16d"0"),(16d"64775"),(16d"64584"),(16d"64936"),(16d"0"),(16d"485"),(16d"621"),(16d"399"),(16d"0"),(16d"65205"),(16d"65109"),(16d"65261"),(16d"0"),(16d"230"),(16d"297"),(16d"192"),(16d"0"),(16d"65377"),(16d"65331"),(16d"65404"),(16d"0"),(16d"108"),(16d"138"),(16d"88"),(16d"0"),(16d"65465"),(16d"65446"),(16d"65479"),(16d"0"),(16d"45"),(16d"56"),(16d"35"),(16d"0"),(16d"65509"),(16d"65502"),(16d"65515"),(16d"0"),(16d"17"),(16d"21"),(16d"14"),(16d"0"),(16d"65524"),(16d"65519"))

	;
end architecture;